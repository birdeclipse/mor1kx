module MEM2_128X16 ( /*AUTOARG*/
   // Outputs
   Q1, Q2,
   // Inputs
   CK1, CK2, CE1, CE2, A1, A2, WE1, WE2, D1, D2
   );

   input CK1;
   input CK2;
   input CE1;
   input CE2;
   input [11:0] A1;
   input [11:0] A2;
   input       WE1;
   input       WE2;
   input [31:0] D1;
   input [31:0] D2;

   output [31:0] Q1;
   output [31:0] Q2;

endmodule
